/home/ykhuang/research/PvsLVS/CurrentMirror_ST/netlist