/home/ykhuang/research/PvsLVS/CurrentSource_All_ST/netlist