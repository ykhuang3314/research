
wire \vdd3! ;

wire \vdde! ;

wire \vdd! ;

wire \gnd! ;
