/home/ykhuang/research/PvsLVS/MultiChannel_ST/netlist