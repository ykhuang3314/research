
wire \gnd! ;

wire \vdd3! ;

wire \vdde! ;

wire \vdd! ;
