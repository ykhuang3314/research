
wire \gnd! ;

wire \vdde! ;

wire \vdd3! ;
