/home/ykhuang/research/PvsLVS/CurrentMirror_x10_LV/netlist