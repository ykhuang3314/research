
wire \gnd! ;
