/home/ykhuang/research/PvsLVS/Ext_Iref_ST/netlist