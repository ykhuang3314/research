/home/ykhuang/research/PvsLVS/Idac_5bit_ST_V2/netlist