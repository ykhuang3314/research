
wire \vdd3! ;

wire \vdde! ;

wire \gnd! ;

wire \vdd! ;
