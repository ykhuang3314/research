
wire \vdd3! ;

wire \vdde! ;

wire \gnd! ;
